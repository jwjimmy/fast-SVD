module scope(clk,a,b,Cout);
